// TestSPI.v

// Generated using ACDS version 11.1sp1 216 at 2012.04.14.18:16:36

`timescale 1 ps / 1 ps
module TestSPI (
		input  wire  reset_reset_n, // reset.reset_n
		input  wire  clk_clk        //   clk.clk
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> spi_0:reset_n

	TestSPI_spi_0 spi_0 (
		.clk           (clk_clk),                         //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset), //            reset.reset_n
		.data_from_cpu (),                                // spi_control_port.writedata
		.data_to_cpu   (),                                //                 .readdata
		.mem_addr      (),                                //                 .address
		.read_n        (),                                //                 .read_n
		.spi_select    (),                                //                 .chipselect
		.write_n       (),                                //                 .write_n
		.dataavailable (),                                //                 .dataavailable
		.endofpacket   (),                                //                 .endofpacket
		.readyfordata  (),                                //                 .readyfordata
		.irq           (),                                //              irq.irq
		.MISO          (),                                //         external.export
		.MOSI          (),                                //                 .export
		.SCLK          (),                                //                 .export
		.SS_n          ()                                 //                 .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
