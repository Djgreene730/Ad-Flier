--	=	=	=	=	=	=	=	=	=	=	=	=	=	=	=
--	Title:		SPI Slave Module
--	Project:	The Ad-Flier, Spring 2012
--	Author:		David Greene
--	=	=	=	=	=	=	=	=	=	=	=	=	=	=	=

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity SPI_Slave is
	port( 
		clk		:	in		std_logic;
		SCK		:	in		std_logic;
		MOSI	:	in		std_logic;
		MISO	:	out		std_logic;
		SSEL	:	in		std_logic;
		LED		:	out		std_logic
	);
end SPI_Slave;

architecture BHV of SPI_Slave is
	
	-- Signals
	signal SCK_risingedge		:	std_logic 						:= '0';
	signal SCK_fallingedge		:	std_logic 						:= '0';
	signal SSEL_active			:	std_logic 						:= '0';
	signal SSEL_startmessage	:	std_logic 						:= '0';
	signal SSEL_endmessage		:	std_logic 						:= '0';
	signal MOSI_data			:	std_logic 						:= '0';
	signal byte_received		:	std_logic 						:= '0';
	signal SCKr					:	std_logic_vector(2 downto 0)	:= (others => '0');
	signal SSELr				:	std_logic_vector(2 downto 0)	:= (others => '0');
	signal MOSIr				:	std_logic_vector(1 downto 0)	:= (others => '0');
	signal bitcnt				:	std_logic_vector(2 downto 0)	:= (others => '0');
	signal byte_data_received	:	std_logic_vector(7 downto 0)	:= (others => '0');
	signal byte_data_sent		:	std_logic_vector(7 downto 0)	:= (others => '0');
	signal cnt					:	std_logic_vector(7 downto 0)	:= (others => '0');

begin
	
	-- Update Registers
	SCK_risingedge		<= '1' when SCKr(2 downto 1) = "01" else '0';		-- Detect SCK Rising Edge
	SCK_fallingedge 	<= '1' when SCKr(2 downto 1) = "10" else '0';		-- Detect SCK Falling Edge
	SSEL_startmessage 	<= '1' when SSELr(2 downto 1) = "10" else '0';	-- Message Starts at Falling Edge of SCK
	SSEL_endmessage 	<= '1' when SSELr(2 downto 1) = "01" else '0';	-- Message Stops at Rising Edge of SCK
	SSEL_active 		<= not SSELr(1);  									-- Select Line is Active Low
	MOSI_data 			<= MOSIr(1);
	
	-- Update SCK Clocks and Counters
	process(clk, SCK, SSEL, MOSI, SCKr, SSELr, MOSIr)
	begin
		if (clk'event and clk = '1') then
			-- Set Simple Signals
			SCKr 	<= 	SCKr(1 downto 0) & SCK;
			SSELr	<=	SSELr(1 downto 0) & SSEL;
			MOSIr	<=	MOSIr(0) & MOSI;

			if (bitcnt = "111") then
				byte_received <= SSEL_active and SCK_risingedge;
			else
				byte_received <= '0';
			end if;
			
			if (byte_received = '1') then
				LED <= byte_data_received(0);
			end if;
			
			if (SSEL_startmessage = '1') then
				cnt <= std_logic_vector(unsigned(cnt) + "00000001");
			end if;
			
		end if;
	end process;

	-- Update Bit_Count & Received-Data Shift Register
	process(clk, SSEL_active, SCK_risingedge, bitcnt, byte_data_received, MOSI_data)
	begin
		if (clk'event and clk = '1') then
			if (SSEL_active = '0') then
				bitcnt <= "000";
			else
				if (SCK_risingedge = '1') then 
					bitcnt <= std_logic_vector(unsigned(bitcnt) + "001");
					byte_data_received <= (byte_data_received(6 downto 0) & MOSI_data);
				end if;
			end if;
		end if;
	end process;


	-- Update Serial Output
	process(clk, SSEL_active, SSEL_startmessage, cnt, SCK_fallingedge, bitcnt, byte_data_sent)
	begin
		if (clk'event and clk = '1') then
			if (SSEL_active = '1') then
				if (SSEL_startmessage = '1') then
					byte_data_sent <= cnt;
				else
					if (SCK_fallingedge = '1') then
						if (bitcnt = "000") then
							byte_data_sent <= (others => '0');
						else
							byte_data_sent <= (byte_data_sent(6 downto 0) & '0');
						end if;
					end if;
				end if;
			end if;
			
			-- Output Highest Bit to Output Line
			MISO <= byte_data_sent(7);			
		end if;
	end process;
	
end BHV; 